`ifndef RAL_USER_REG_MODEL_PKG
`define RAL_USER_REG_MODEL_PKG

package ral_user_reg_model_pkg;
import uvm_pkg::*;

class ral_reg_user_reg_model_GDMA_MISC_CONF_REG extends uvm_reg;
	uvm_reg_field resvered1;
	rand uvm_reg_field gdma_ahbm_rst_inter;
	rand uvm_reg_field gdma_arb_pri_dis;
	uvm_reg_field resvered0;
	rand uvm_reg_field gdma_clk_en;
   local uvm_reg_data_t m_data;
   local uvm_reg_data_t m_be;
   local bit            m_is_read;

	covergroup cg_bits ();
	   option.per_instance = 1;
	   option.name = get_name();
	   resvered1: coverpoint {m_data[31:4], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {29'b???????????????????????????00};
	      wildcard bins bit_0_wr_as_1 = {29'b???????????????????????????10};
	      wildcard bins bit_0_rd = {29'b????????????????????????????1};
	      wildcard bins bit_1_wr_as_0 = {29'b??????????????????????????0?0};
	      wildcard bins bit_1_wr_as_1 = {29'b??????????????????????????1?0};
	      wildcard bins bit_1_rd = {29'b????????????????????????????1};
	      wildcard bins bit_2_wr_as_0 = {29'b?????????????????????????0??0};
	      wildcard bins bit_2_wr_as_1 = {29'b?????????????????????????1??0};
	      wildcard bins bit_2_rd = {29'b????????????????????????????1};
	      wildcard bins bit_3_wr_as_0 = {29'b????????????????????????0???0};
	      wildcard bins bit_3_wr_as_1 = {29'b????????????????????????1???0};
	      wildcard bins bit_3_rd = {29'b????????????????????????????1};
	      wildcard bins bit_4_wr_as_0 = {29'b???????????????????????0????0};
	      wildcard bins bit_4_wr_as_1 = {29'b???????????????????????1????0};
	      wildcard bins bit_4_rd = {29'b????????????????????????????1};
	      wildcard bins bit_5_wr_as_0 = {29'b??????????????????????0?????0};
	      wildcard bins bit_5_wr_as_1 = {29'b??????????????????????1?????0};
	      wildcard bins bit_5_rd = {29'b????????????????????????????1};
	      wildcard bins bit_6_wr_as_0 = {29'b?????????????????????0??????0};
	      wildcard bins bit_6_wr_as_1 = {29'b?????????????????????1??????0};
	      wildcard bins bit_6_rd = {29'b????????????????????????????1};
	      wildcard bins bit_7_wr_as_0 = {29'b????????????????????0???????0};
	      wildcard bins bit_7_wr_as_1 = {29'b????????????????????1???????0};
	      wildcard bins bit_7_rd = {29'b????????????????????????????1};
	      wildcard bins bit_8_wr_as_0 = {29'b???????????????????0????????0};
	      wildcard bins bit_8_wr_as_1 = {29'b???????????????????1????????0};
	      wildcard bins bit_8_rd = {29'b????????????????????????????1};
	      wildcard bins bit_9_wr_as_0 = {29'b??????????????????0?????????0};
	      wildcard bins bit_9_wr_as_1 = {29'b??????????????????1?????????0};
	      wildcard bins bit_9_rd = {29'b????????????????????????????1};
	      wildcard bins bit_10_wr_as_0 = {29'b?????????????????0??????????0};
	      wildcard bins bit_10_wr_as_1 = {29'b?????????????????1??????????0};
	      wildcard bins bit_10_rd = {29'b????????????????????????????1};
	      wildcard bins bit_11_wr_as_0 = {29'b????????????????0???????????0};
	      wildcard bins bit_11_wr_as_1 = {29'b????????????????1???????????0};
	      wildcard bins bit_11_rd = {29'b????????????????????????????1};
	      wildcard bins bit_12_wr_as_0 = {29'b???????????????0????????????0};
	      wildcard bins bit_12_wr_as_1 = {29'b???????????????1????????????0};
	      wildcard bins bit_12_rd = {29'b????????????????????????????1};
	      wildcard bins bit_13_wr_as_0 = {29'b??????????????0?????????????0};
	      wildcard bins bit_13_wr_as_1 = {29'b??????????????1?????????????0};
	      wildcard bins bit_13_rd = {29'b????????????????????????????1};
	      wildcard bins bit_14_wr_as_0 = {29'b?????????????0??????????????0};
	      wildcard bins bit_14_wr_as_1 = {29'b?????????????1??????????????0};
	      wildcard bins bit_14_rd = {29'b????????????????????????????1};
	      wildcard bins bit_15_wr_as_0 = {29'b????????????0???????????????0};
	      wildcard bins bit_15_wr_as_1 = {29'b????????????1???????????????0};
	      wildcard bins bit_15_rd = {29'b????????????????????????????1};
	      wildcard bins bit_16_wr_as_0 = {29'b???????????0????????????????0};
	      wildcard bins bit_16_wr_as_1 = {29'b???????????1????????????????0};
	      wildcard bins bit_16_rd = {29'b????????????????????????????1};
	      wildcard bins bit_17_wr_as_0 = {29'b??????????0?????????????????0};
	      wildcard bins bit_17_wr_as_1 = {29'b??????????1?????????????????0};
	      wildcard bins bit_17_rd = {29'b????????????????????????????1};
	      wildcard bins bit_18_wr_as_0 = {29'b?????????0??????????????????0};
	      wildcard bins bit_18_wr_as_1 = {29'b?????????1??????????????????0};
	      wildcard bins bit_18_rd = {29'b????????????????????????????1};
	      wildcard bins bit_19_wr_as_0 = {29'b????????0???????????????????0};
	      wildcard bins bit_19_wr_as_1 = {29'b????????1???????????????????0};
	      wildcard bins bit_19_rd = {29'b????????????????????????????1};
	      wildcard bins bit_20_wr_as_0 = {29'b???????0????????????????????0};
	      wildcard bins bit_20_wr_as_1 = {29'b???????1????????????????????0};
	      wildcard bins bit_20_rd = {29'b????????????????????????????1};
	      wildcard bins bit_21_wr_as_0 = {29'b??????0?????????????????????0};
	      wildcard bins bit_21_wr_as_1 = {29'b??????1?????????????????????0};
	      wildcard bins bit_21_rd = {29'b????????????????????????????1};
	      wildcard bins bit_22_wr_as_0 = {29'b?????0??????????????????????0};
	      wildcard bins bit_22_wr_as_1 = {29'b?????1??????????????????????0};
	      wildcard bins bit_22_rd = {29'b????????????????????????????1};
	      wildcard bins bit_23_wr_as_0 = {29'b????0???????????????????????0};
	      wildcard bins bit_23_wr_as_1 = {29'b????1???????????????????????0};
	      wildcard bins bit_23_rd = {29'b????????????????????????????1};
	      wildcard bins bit_24_wr_as_0 = {29'b???0????????????????????????0};
	      wildcard bins bit_24_wr_as_1 = {29'b???1????????????????????????0};
	      wildcard bins bit_24_rd = {29'b????????????????????????????1};
	      wildcard bins bit_25_wr_as_0 = {29'b??0?????????????????????????0};
	      wildcard bins bit_25_wr_as_1 = {29'b??1?????????????????????????0};
	      wildcard bins bit_25_rd = {29'b????????????????????????????1};
	      wildcard bins bit_26_wr_as_0 = {29'b?0??????????????????????????0};
	      wildcard bins bit_26_wr_as_1 = {29'b?1??????????????????????????0};
	      wildcard bins bit_26_rd = {29'b????????????????????????????1};
	      wildcard bins bit_27_wr_as_0 = {29'b0???????????????????????????0};
	      wildcard bins bit_27_wr_as_1 = {29'b1???????????????????????????0};
	      wildcard bins bit_27_rd = {29'b????????????????????????????1};
	      option.weight = 84;
	   }
	   gdma_ahbm_rst_inter: coverpoint {m_data[3:3], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   gdma_arb_pri_dis: coverpoint {m_data[2:2], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	   resvered0: coverpoint {m_data[1:1], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd = {2'b?1};
	      option.weight = 3;
	   }
	   gdma_clk_en: coverpoint {m_data[0:0], m_is_read} iff(m_be) {
	      wildcard bins bit_0_wr_as_0 = {2'b00};
	      wildcard bins bit_0_wr_as_1 = {2'b10};
	      wildcard bins bit_0_rd_as_0 = {2'b01};
	      wildcard bins bit_0_rd_as_1 = {2'b11};
	      option.weight = 4;
	   }
	endgroup
	covergroup cg_vals ();
		option.per_instance = 1;
		resvered1_value : coverpoint resvered1.value {
			bins min = { 28'h0 };
			bins max = { 28'hFFFFFFF };
			bins others = { [28'h1:28'hFFFFFFE] };
			option.weight = 3;
		}
		gdma_ahbm_rst_inter_value : coverpoint gdma_ahbm_rst_inter.value[0:0] {
			option.weight = 2;
		}
		gdma_arb_pri_dis_value : coverpoint gdma_arb_pri_dis.value[0:0] {
			option.weight = 2;
		}
		resvered0_value : coverpoint resvered0.value[0:0] {
			option.weight = 2;
		}
		gdma_clk_en_value : coverpoint gdma_clk_en.value[0:0] {
			option.weight = 2;
		}
	endgroup : cg_vals

	function new(string name = "user_reg_model_GDMA_MISC_CONF_REG");
		super.new(name, 32,build_coverage(UVM_CVR_REG_BITS+UVM_CVR_FIELD_VALS));
		if (has_coverage(UVM_CVR_REG_BITS))
			cg_bits = new();
		if (has_coverage(UVM_CVR_FIELD_VALS))
			cg_vals = new();
	endfunction: new
   virtual function void build();
      this.resvered1 = uvm_reg_field::type_id::create("resvered1",,get_full_name());
      this.resvered1.configure(this, 28, 4, "RO", 0, 28'b0, 1, 0, 0);
      this.gdma_ahbm_rst_inter = uvm_reg_field::type_id::create("gdma_ahbm_rst_inter",,get_full_name());
      this.gdma_ahbm_rst_inter.configure(this, 1, 3, "RW", 0, 1'b1, 1, 0, 0);
      this.gdma_arb_pri_dis = uvm_reg_field::type_id::create("gdma_arb_pri_dis",,get_full_name());
      this.gdma_arb_pri_dis.configure(this, 1, 2, "RW", 0, 1'b0, 1, 0, 0);
      this.resvered0 = uvm_reg_field::type_id::create("resvered0",,get_full_name());
      this.resvered0.configure(this, 1, 1, "RO", 0, 1'b0, 1, 0, 0);
      this.gdma_clk_en = uvm_reg_field::type_id::create("gdma_clk_en",,get_full_name());
      this.gdma_clk_en.configure(this, 1, 0, "RW", 0, 1'b1, 1, 0, 0);
   endfunction: build

	`uvm_object_utils(ral_reg_user_reg_model_GDMA_MISC_CONF_REG)


	virtual function void sample(uvm_reg_data_t data,
	                             uvm_reg_data_t byte_en,
	                             bit            is_read,
	                             uvm_reg_map    map);
	   if (get_coverage(UVM_CVR_REG_BITS)) begin
	      m_data    = data;
	      m_be      = byte_en;
	      m_is_read = is_read;
	      cg_bits.sample();
	   end
	endfunction

	function void sample_values();
	   super.sample_values();
	   if (get_coverage(UVM_CVR_FIELD_VALS)) begin
	      if(cg_vals!=null) cg_vals.sample();
	   end
	endfunction
endclass : ral_reg_user_reg_model_GDMA_MISC_CONF_REG


class ral_mem_user_reg_model_tx_ram extends uvm_mem;
   function new(string name = "user_reg_model_tx_ram");
      super.new(name, `UVM_REG_ADDR_WIDTH'h20, 128, "RW", build_coverage(UVM_CVR_ADDR_MAP));
   endfunction
   virtual function void build();
   endfunction: build

   `uvm_object_utils(ral_mem_user_reg_model_tx_ram)

endclass : ral_mem_user_reg_model_tx_ram


class ral_block_user_reg_model extends uvm_reg_block;
	rand ral_reg_user_reg_model_GDMA_MISC_CONF_REG GDMA_MISC_CONF_REG;
	rand ral_mem_user_reg_model_tx_ram tx_ram;
   local uvm_reg_data_t m_offset;
	uvm_reg_field GDMA_MISC_CONF_REG_resvered1;
	uvm_reg_field resvered1;
	rand uvm_reg_field GDMA_MISC_CONF_REG_gdma_ahbm_rst_inter;
	rand uvm_reg_field gdma_ahbm_rst_inter;
	rand uvm_reg_field GDMA_MISC_CONF_REG_gdma_arb_pri_dis;
	rand uvm_reg_field gdma_arb_pri_dis;
	uvm_reg_field GDMA_MISC_CONF_REG_resvered0;
	uvm_reg_field resvered0;
	rand uvm_reg_field GDMA_MISC_CONF_REG_gdma_clk_en;
	rand uvm_reg_field gdma_clk_en;


covergroup cg_addr (input string name);
	option.per_instance = 1;
option.name = get_name();

	GDMA_MISC_CONF_REG : coverpoint m_offset {
		bins accessed = { `UVM_REG_ADDR_WIDTH'h44 };
		option.weight = 1;
	}

	tx_ram : coverpoint m_offset {
		bins first_location_accessed = { [`UVM_REG_ADDR_WIDTH'hFF:`UVM_REG_ADDR_WIDTH'h102] };
		bins last_location_accessed = { [`UVM_REG_ADDR_WIDTH'h17B:`UVM_REG_ADDR_WIDTH'h17E] };
		bins other_locations_accessed = { [`UVM_REG_ADDR_WIDTH'h103:`UVM_REG_ADDR_WIDTH'h17A] };
		option.weight = 3;
	}
endgroup
	function new(string name = "user_reg_model");
		super.new(name, build_coverage(UVM_CVR_ADDR_MAP+UVM_CVR_FIELD_VALS));
		if (has_coverage(UVM_CVR_ADDR_MAP))
			cg_addr = new("cg_addr");
	endfunction: new

   virtual function void build();
      this.default_map = create_map("", 0, 4, UVM_LITTLE_ENDIAN, 0);
      this.GDMA_MISC_CONF_REG = ral_reg_user_reg_model_GDMA_MISC_CONF_REG::type_id::create("GDMA_MISC_CONF_REG",,get_full_name());
      if(this.GDMA_MISC_CONF_REG.has_coverage(UVM_CVR_REG_BITS))
      	this.GDMA_MISC_CONF_REG.cg_bits.option.name = {get_name(), ".", "GDMA_MISC_CONF_REG_bits"};
      this.GDMA_MISC_CONF_REG.configure(this, null, "");
      this.GDMA_MISC_CONF_REG.build();
         this.GDMA_MISC_CONF_REG.add_hdl_path('{
            '{"resvered1", 4, 28},
            '{"gdma_ahbm_rst_inter", 3, 1},
            '{"gdma_arb_pri_dis", 2, 1},
            '{"resvered0", 1, 1},
            '{"gdma_clk_en", 0, 1}
         });
      this.default_map.add_reg(this.GDMA_MISC_CONF_REG, `UVM_REG_ADDR_WIDTH'h44, "RW", 0);
		this.GDMA_MISC_CONF_REG_resvered1 = this.GDMA_MISC_CONF_REG.resvered1;
		this.resvered1 = this.GDMA_MISC_CONF_REG.resvered1;
		this.GDMA_MISC_CONF_REG_gdma_ahbm_rst_inter = this.GDMA_MISC_CONF_REG.gdma_ahbm_rst_inter;
		this.gdma_ahbm_rst_inter = this.GDMA_MISC_CONF_REG.gdma_ahbm_rst_inter;
		this.GDMA_MISC_CONF_REG_gdma_arb_pri_dis = this.GDMA_MISC_CONF_REG.gdma_arb_pri_dis;
		this.gdma_arb_pri_dis = this.GDMA_MISC_CONF_REG.gdma_arb_pri_dis;
		this.GDMA_MISC_CONF_REG_resvered0 = this.GDMA_MISC_CONF_REG.resvered0;
		this.resvered0 = this.GDMA_MISC_CONF_REG.resvered0;
		this.GDMA_MISC_CONF_REG_gdma_clk_en = this.GDMA_MISC_CONF_REG.gdma_clk_en;
		this.gdma_clk_en = this.GDMA_MISC_CONF_REG.gdma_clk_en;
      this.tx_ram = ral_mem_user_reg_model_tx_ram::type_id::create("tx_ram",,get_full_name());
      this.tx_ram.configure(this, "");
      this.tx_ram.build();
      this.default_map.add_mem(this.tx_ram, `UVM_REG_ADDR_WIDTH'hFF, "RW", 0);
   endfunction : build

	`uvm_object_utils(ral_block_user_reg_model)


function void sample(uvm_reg_addr_t offset,
                     bit            is_read,
                     uvm_reg_map    map);
  if (get_coverage(UVM_CVR_ADDR_MAP)) begin
    m_offset = offset;
    cg_addr.sample();
  end
endfunction

	function void sample_values();
	   super.sample_values();
		if (get_coverage(UVM_CVR_FIELD_VALS)) begin
			if (GDMA_MISC_CONF_REG.cg_vals != null) GDMA_MISC_CONF_REG.cg_vals.sample();
		end
	endfunction
endclass : ral_block_user_reg_model


endpackage
`endif
